module debounce_input
#(
)
(
);



endmodule
