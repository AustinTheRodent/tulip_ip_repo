module half_band_brom
(
  input  logic        clk,

  input  logic [7:0]  din_address,
  input  logic        din_valid,

  output logic [15:0] dout,
  output logic        dout_valid
);

  logic signed [15:0] brom_data [0:2**8-1] =
  {
    25            ,
    -54           ,
    -26           ,
    2             ,
    8             ,
    -10           ,
    -12           ,
    9             ,
    14            ,
    -9            ,
    -16           ,
    9             ,
    17            ,
    -9            ,
    -20           ,
    8             ,
    22            ,
    -7            ,
    -24           ,
    6             ,
    26            ,
    -5            ,
    -29           ,
    4             ,
    31            ,
    -2            ,
    -34           ,
    0             ,
    36            ,
    2             ,
    -39           ,
    -5            ,
    41            ,
    8             ,
    -43           ,
    -11           ,
    46            ,
    15            ,
    -48           ,
    -19           ,
    50            ,
    24            ,
    -51           ,
    -29           ,
    53            ,
    34            ,
    -54           ,
    -40           ,
    55            ,
    46            ,
    -55           ,
    -52           ,
    55            ,
    59            ,
    -55           ,
    -66           ,
    54            ,
    73            ,
    -52           ,
    -81           ,
    50            ,
    89            ,
    -48           ,
    -98           ,
    44            ,
    107           ,
    -40           ,
    -116          ,
    35            ,
    125           ,
    -29           ,
    -134          ,
    22            ,
    144           ,
    -14           ,
    -154          ,
    5             ,
    163           ,
    5             ,
    -173          ,
    -17           ,
    183           ,
    30            ,
    -193          ,
    -44           ,
    203           ,
    60            ,
    -213          ,
    -78           ,
    222           ,
    98            ,
    -232          ,
    -120          ,
    241           ,
    145           ,
    -250          ,
    -173          ,
    259           ,
    204           ,
    -267          ,
    -239          ,
    275           ,
    279           ,
    -282          ,
    -324          ,
    289           ,
    377           ,
    -296          ,
    -440          ,
    302           ,
    515           ,
    -307          ,
    -608          ,
    312           ,
    727           ,
    -317          ,
    -885          ,
    320           ,
    1108          ,
    -323          ,
    -1452         ,
    326           ,
    2063          ,
    -327          ,
    -3471         ,
    328           ,
    10461         ,
    16113         ,
    10461         ,
    328           ,
    -3471         ,
    -327          ,
    2063          ,
    326           ,
    -1452         ,
    -323          ,
    1108          ,
    320           ,
    -885          ,
    -317          ,
    727           ,
    312           ,
    -608          ,
    -307          ,
    515           ,
    302           ,
    -440          ,
    -296          ,
    377           ,
    289           ,
    -324          ,
    -282          ,
    279           ,
    275           ,
    -239          ,
    -267          ,
    204           ,
    259           ,
    -173          ,
    -250          ,
    145           ,
    241           ,
    -120          ,
    -232          ,
    98            ,
    222           ,
    -78           ,
    -213          ,
    60            ,
    203           ,
    -44           ,
    -193          ,
    30            ,
    183           ,
    -17           ,
    -173          ,
    5             ,
    163           ,
    5             ,
    -154          ,
    -14           ,
    144           ,
    22            ,
    -134          ,
    -29           ,
    125           ,
    35            ,
    -116          ,
    -40           ,
    107           ,
    44            ,
    -98           ,
    -48           ,
    89            ,
    50            ,
    -81           ,
    -52           ,
    73            ,
    54            ,
    -66           ,
    -55           ,
    59            ,
    55            ,
    -52           ,
    -55           ,
    46            ,
    55            ,
    -40           ,
    -54           ,
    34            ,
    53            ,
    -29           ,
    -51           ,
    24            ,
    50            ,
    -19           ,
    -48           ,
    15            ,
    46            ,
    -11           ,
    -43           ,
    8             ,
    41            ,
    -5            ,
    -39           ,
    2             ,
    36            ,
    0             ,
    -34           ,
    -2            ,
    31            ,
    4             ,
    -29           ,
    -5            ,
    26            ,
    6             ,
    -24           ,
    -7            ,
    22            ,
    8             ,
    -20           ,
    -9            ,
    17            ,
    9             ,
    -16           ,
    -9            ,
    14            ,
    9             ,
    -12           ,
    -10           ,
    8             ,
    2             ,
    -26           ,
    -54           ,
    25            ,
    0
  };

/////////////////////////////////////////////////////////////////////

  always @ (posedge clk) begin
    dout        <= brom_data[din_address];
    dout_valid  <= din_valid;
  end

endmodule
