module half_band_brom
(
  input  logic        clk,

  input  logic [8:0]  din_address,
  input  logic        din_valid,

  output logic [15:0] dout,
  output logic        dout_valid
);

  logic signed [15:0] brom_data [0:2**9-1] =
  {
    61               ,
    113              ,
    -54              ,
    13               ,
    -1               ,
    11               ,
    -9               ,
    -7               ,
    7                ,
    8                ,
    -8               ,
    -9               ,
    8                ,
    9                ,
    -8               ,
    -10              ,
    8                ,
    10               ,
    -8               ,
    -11              ,
    8                ,
    11               ,
    -8               ,
    -12              ,
    8                ,
    12               ,
    -8               ,
    -13              ,
    8                ,
    13               ,
    -8               ,
    -14              ,
    8                ,
    15               ,
    -8               ,
    -15              ,
    8                ,
    16               ,
    -8               ,
    -16              ,
    8                ,
    17               ,
    -8               ,
    -18              ,
    8                ,
    18               ,
    -8               ,
    -19              ,
    8                ,
    20               ,
    -8               ,
    -21              ,
    7                ,
    21               ,
    -7               ,
    -22              ,
    7                ,
    23               ,
    -7               ,
    -24              ,
    7                ,
    24               ,
    -6               ,
    -25              ,
    6                ,
    26               ,
    -6               ,
    -27              ,
    5                ,
    28               ,
    -5               ,
    -28              ,
    4                ,
    29               ,
    -4               ,
    -30              ,
    4                ,
    31               ,
    -3               ,
    -32              ,
    3                ,
    33               ,
    -2               ,
    -34              ,
    1                ,
    35               ,
    -1               ,
    -36              ,
    0                ,
    37               ,
    1                ,
    -38              ,
    -1               ,
    38               ,
    2                ,
    -39              ,
    -3               ,
    40               ,
    4                ,
    -41              ,
    -5               ,
    42               ,
    6                ,
    -43              ,
    -7               ,
    44               ,
    8                ,
    -45              ,
    -9               ,
    46               ,
    10               ,
    -47              ,
    -11              ,
    48               ,
    12               ,
    -49              ,
    -13              ,
    50               ,
    15               ,
    -51              ,
    -16              ,
    52               ,
    17               ,
    -53              ,
    -19              ,
    54               ,
    20               ,
    -56              ,
    -22              ,
    57               ,
    24               ,
    -58              ,
    -25              ,
    59               ,
    27               ,
    -60              ,
    -29              ,
    61               ,
    31               ,
    -62              ,
    -33              ,
    63               ,
    35               ,
    -64              ,
    -37              ,
    65               ,
    39               ,
    -66              ,
    -42              ,
    67               ,
    44               ,
    -68              ,
    -47              ,
    69               ,
    49               ,
    -70              ,
    -52              ,
    71               ,
    55               ,
    -72              ,
    -58              ,
    72               ,
    61               ,
    -73              ,
    -64              ,
    74               ,
    67               ,
    -75              ,
    -71              ,
    76               ,
    74               ,
    -77              ,
    -78              ,
    78               ,
    82               ,
    -79              ,
    -86              ,
    80               ,
    90               ,
    -80              ,
    -95              ,
    81               ,
    99               ,
    -82              ,
    -104             ,
    83               ,
    109              ,
    -84              ,
    -115             ,
    84               ,
    121              ,
    -85              ,
    -127             ,
    86               ,
    133              ,
    -87              ,
    -140             ,
    87               ,
    147              ,
    -88              ,
    -155             ,
    89               ,
    163              ,
    -89              ,
    -172             ,
    90               ,
    181              ,
    -90              ,
    -191             ,
    91               ,
    202              ,
    -91              ,
    -214             ,
    92               ,
    227              ,
    -92              ,
    -241             ,
    93               ,
    256              ,
    -93              ,
    -274             ,
    94               ,
    293              ,
    -94              ,
    -314             ,
    95               ,
    338              ,
    -95              ,
    -366             ,
    95               ,
    398              ,
    -96              ,
    -435             ,
    96               ,
    479              ,
    -96              ,
    -532             ,
    96               ,
    598              ,
    -97              ,
    -680             ,
    97               ,
    787              ,
    -97              ,
    -933             ,
    97               ,
    1144             ,
    -97              ,
    -1473            ,
    97               ,
    2066             ,
    -97              ,
    -3446            ,
    97               ,
    10344            ,
    16152            ,
    10344            ,
    97               ,
    -3446            ,
    -97              ,
    2066             ,
    97               ,
    -1473            ,
    -97              ,
    1144             ,
    97               ,
    -933             ,
    -97              ,
    787              ,
    97               ,
    -680             ,
    -97              ,
    598              ,
    96               ,
    -532             ,
    -96              ,
    479              ,
    96               ,
    -435             ,
    -96              ,
    398              ,
    95               ,
    -366             ,
    -95              ,
    338              ,
    95               ,
    -314             ,
    -94              ,
    293              ,
    94               ,
    -274             ,
    -93              ,
    256              ,
    93               ,
    -241             ,
    -92              ,
    227              ,
    92               ,
    -214             ,
    -91              ,
    202              ,
    91               ,
    -191             ,
    -90              ,
    181              ,
    90               ,
    -172             ,
    -89              ,
    163              ,
    89               ,
    -155             ,
    -88              ,
    147              ,
    87               ,
    -140             ,
    -87              ,
    133              ,
    86               ,
    -127             ,
    -85              ,
    121              ,
    84               ,
    -115             ,
    -84              ,
    109              ,
    83               ,
    -104             ,
    -82              ,
    99               ,
    81               ,
    -95              ,
    -80              ,
    90               ,
    80               ,
    -86              ,
    -79              ,
    82               ,
    78               ,
    -78              ,
    -77              ,
    74               ,
    76               ,
    -71              ,
    -75              ,
    67               ,
    74               ,
    -64              ,
    -73              ,
    61               ,
    72               ,
    -58              ,
    -72              ,
    55               ,
    71               ,
    -52              ,
    -70              ,
    49               ,
    69               ,
    -47              ,
    -68              ,
    44               ,
    67               ,
    -42              ,
    -66              ,
    39               ,
    65               ,
    -37              ,
    -64              ,
    35               ,
    63               ,
    -33              ,
    -62              ,
    31               ,
    61               ,
    -29              ,
    -60              ,
    27               ,
    59               ,
    -25              ,
    -58              ,
    24               ,
    57               ,
    -22              ,
    -56              ,
    20               ,
    54               ,
    -19              ,
    -53              ,
    17               ,
    52               ,
    -16              ,
    -51              ,
    15               ,
    50               ,
    -13              ,
    -49              ,
    12               ,
    48               ,
    -11              ,
    -47              ,
    10               ,
    46               ,
    -9               ,
    -45              ,
    8                ,
    44               ,
    -7               ,
    -43              ,
    6                ,
    42               ,
    -5               ,
    -41              ,
    4                ,
    40               ,
    -3               ,
    -39              ,
    2                ,
    38               ,
    -1               ,
    -38              ,
    1                ,
    37               ,
    0                ,
    -36              ,
    -1               ,
    35               ,
    1                ,
    -34              ,
    -2               ,
    33               ,
    3                ,
    -32              ,
    -3               ,
    31               ,
    4                ,
    -30              ,
    -4               ,
    29               ,
    4                ,
    -28              ,
    -5               ,
    28               ,
    5                ,
    -27              ,
    -6               ,
    26               ,
    6                ,
    -25              ,
    -6               ,
    24               ,
    7                ,
    -24              ,
    -7               ,
    23               ,
    7                ,
    -22              ,
    -7               ,
    21               ,
    7                ,
    -21              ,
    -8               ,
    20               ,
    8                ,
    -19              ,
    -8               ,
    18               ,
    8                ,
    -18              ,
    -8               ,
    17               ,
    8                ,
    -16              ,
    -8               ,
    16               ,
    8                ,
    -15              ,
    -8               ,
    15               ,
    8                ,
    -14              ,
    -8               ,
    13               ,
    8                ,
    -13              ,
    -8               ,
    12               ,
    8                ,
    -12              ,
    -8               ,
    11               ,
    8                ,
    -11              ,
    -8               ,
    10               ,
    8                ,
    -10              ,
    -8               ,
    9                ,
    8                ,
    -9               ,
    -8               ,
    8                ,
    7                ,
    -7               ,
    -9               ,
    11               ,
    -1               ,
    13               ,
    -54              ,
    113              ,
    61               ,
    0
  };

/////////////////////////////////////////////////////////////////////

  always @ (posedge clk) begin
    dout        <= brom_data[din_address];
    dout_valid  <= din_valid;
  end

endmodule
